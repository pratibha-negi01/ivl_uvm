..j
